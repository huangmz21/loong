`include "mycpu.h"

module wb_stage(
    input                           clk           ,
    input                           reset         ,
    //allowin
    output                          ws_allowin    ,
    //from ms
    input                           ms_to_ws_valid,
    input  [`MS_TO_WS_BUS_WD -1:0]  ms_to_ws_bus  ,
    //to rf: for write back
    output [`WS_TO_RF_BUS_WD -1:0]  ws_to_rf_bus  ,
    //forwardpath
    output [32-1:0]                 es_forward_ws,
    //trace debug interface
    output [31:0] debug_wb_pc     ,
    output [ 3:0] debug_wb_rf_wen ,
    output [ 4:0] debug_wb_rf_wnum,
    output [31:0] debug_wb_rf_wdata
);

 (* keep = "true" *) reg         ws_valid;
wire        ws_ready_go;

 (* keep = "true" *) reg [`MS_TO_WS_BUS_WD -1:0] ms_to_ws_bus_r;
 //////1
wire        ws_res_from_mem_h;
wire        ws_res_from_mem_b;
wire        ws_res_from_mem_sign;
wire [1:0]  ws_whb_mux;
//////0
wire        ws_gr_we;
wire [ 4:0] ws_dest;
wire [31:0] ws_final_result;
wire [31:0] ws_pc;
assign {//////1
        ws_res_from_mem_h,  //74:74
        ws_res_from_mem_b,  //73:73
        ws_res_from_mem_sign,//72:72
        ws_whb_mux,//71:70
        //////1
        ws_gr_we       ,  //69:69
        ws_dest        ,  //68:64
        ws_final_result,  //63:32
        ws_pc             //31:0
       } = ms_to_ws_bus_r;

wire        rf_we;
wire [4 :0] rf_waddr;
wire [31:0] rf_wdata;
assign ws_to_rf_bus = {rf_we   ,  //37:37
                       rf_waddr,  //36:32
                       rf_wdata   //31:0
                      };

assign ws_ready_go = 1'b1;
assign ws_allowin  = !ws_valid || ws_ready_go;
always @(posedge clk) begin
    if (reset) begin
        ws_valid <= 1'b0;
    end
    else if (ws_allowin) begin
        ws_valid <= ms_to_ws_valid;
    end

    if (ms_to_ws_valid && ws_allowin) begin
        ms_to_ws_bus_r <= ms_to_ws_bus;
    end
end

assign rf_we    = ws_gr_we&&ws_valid;
assign rf_waddr = ws_dest;
assign rf_wdata = (ws_res_from_mem_h && ~ws_whb_mux[1] && ws_res_from_mem_sign) ? {{16{ws_final_result[15]}}, ws_final_result[15:0]} :
                  (ws_res_from_mem_h && ~ws_whb_mux[1] &&~ws_res_from_mem_sign) ? {{16{1'b0}}, ws_final_result[15:0]} :
                  (ws_res_from_mem_h &&  ws_whb_mux[1] && ws_res_from_mem_sign) ? {{16{ws_final_result[31]}}, ws_final_result[31:16]} :
                  (ws_res_from_mem_h &&  ws_whb_mux[1] &&~ws_res_from_mem_sign) ? {{16{1'b0}}, ws_final_result[31:16]} :
                  (ws_res_from_mem_b && ~ws_whb_mux[1] && ~ws_whb_mux[0] && ws_res_from_mem_sign) ? {{24{ws_final_result[7]}}, ws_final_result[7:0]} :
                  (ws_res_from_mem_b && ~ws_whb_mux[1] && ~ws_whb_mux[0] &&~ws_res_from_mem_sign) ? {{24{1'b0}}, ws_final_result[7:0]} :
                  (ws_res_from_mem_b && ~ws_whb_mux[1] &&  ws_whb_mux[0] && ws_res_from_mem_sign) ? {{24{ws_final_result[15]}}, ws_final_result[15:8]} :
                  (ws_res_from_mem_b && ~ws_whb_mux[1] &&  ws_whb_mux[0] &&~ws_res_from_mem_sign) ? {{24{1'b0}}, ws_final_result[15:8]} :
                  (ws_res_from_mem_b &&  ws_whb_mux[1] && ~ws_whb_mux[0] && ws_res_from_mem_sign) ? {{24{ws_final_result[23]}}, ws_final_result[23:16]} :
                  (ws_res_from_mem_b &&  ws_whb_mux[1] && ~ws_whb_mux[0] &&~ws_res_from_mem_sign) ? {{24{1'b0}}, ws_final_result[23:16]} :
                  (ws_res_from_mem_b &&  ws_whb_mux[1] &&  ws_whb_mux[0] && ws_res_from_mem_sign) ? {{24{ws_final_result[31]}}, ws_final_result[31:24]} :
                  (ws_res_from_mem_b &&  ws_whb_mux[1] &&  ws_whb_mux[0] &&~ws_res_from_mem_sign) ? {{24{1'b0}}, ws_final_result[31:24]} :
                   ws_final_result;
assign es_forward_ws = ws_final_result;/////是否改成rf_wdata？

// debug info generate
assign debug_wb_pc       = ws_pc;
assign debug_wb_rf_wen   = {4{rf_we}};
assign debug_wb_rf_wnum  = ws_dest;
//////1
assign debug_wb_rf_wdata = rf_wdata;
//////0

endmodule
